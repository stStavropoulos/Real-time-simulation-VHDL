library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_textio.all;
use std.textio.all;

Package readdatapart1 is
type bk is array (1 to 3) of std_logic_vector(34 downto 0);
type A0 is array (1 to 3,1 to 3) of signed(34 downto 0);
type history1 is array (1 to 2,1 to 4) of signed(34 downto 0);
type history2 is array (1 to 6,1 to 4) of signed(34 downto 0);
type matrix is array (1 to 9) of std_logic_vector(34 downto 0);
type part_mat is array (1 to 200) of std_logic_vector(34 downto 0);
type single is array(1 to 6) of std_logic_vector(34 downto 0);
type values is array(1 to 40) of std_logic_vector(34 downto 0);
impure function readmatrix(constant MatFilename: in string) return matrix; 
impure function readmatrix2 (constant MatFilename : in string) return part_mat ;
impure function readmatrix3 (constant MatFilename : in string) return single ;
impure function readmatrix4 (constant MatFilename : in string) return values ;
end readdatapart1;

Package body readdatapart1 is

impure function readmatrix (constant MatFilename : in string) return matrix is
FILE MatFile : text is in MatFileName;
variable MatFileLine : line;
variable Mat : matrix;
begin
for i in 1 to 9 loop
readline (MatFile, MatFileLine);
read (MatFileLine, Mat(i));
end loop;
return Mat;
end function; 


impure function readmatrix2 (constant MatFilename : in string) return part_mat is
FILE MatFile : text is in MatFileName;
variable MatFileLine : line;
variable Mat_p : part_mat;
begin
for i in 1 to 200 loop
readline (MatFile, MatFileLine);
read (MatFileLine, Mat_p(i));
end loop;
return Mat_p;
end function; 

impure function readmatrix3 (constant MatFilename : in string) return single is
FILE MatFile : text is in MatFileName;
variable MatFileLine : line;
variable Mat_p : single;
begin
for i in 1 to 6 loop
readline (MatFile, MatFileLine);
read (MatFileLine, Mat_p(i));
end loop;
return Mat_p;
end function; 

impure function readmatrix4 (constant MatFilename : in string) return values is
FILE MatFile : text is in MatFileName;
variable MatFileLine : line;
variable Mat_p : values;
begin
for i in 1 to 40 loop
readline (MatFile, MatFileLine);
read (MatFileLine, Mat_p(i));
end loop;
return Mat_p;
end function; 



end readdatapart1;